module matriz_mul_escalar(matrizA, scl, matriz_resultante);
	input [199:0] matrizA;
	input [7:0] scl;
	output wire [199:0] matriz_resultante;
	
	genvar i;
	
	generate
		for (i = 0; i < 25; i = i + 1) begin : soma_matrizes
			assign matriz_resultante[i*8 +: 8] = scl * matrizA[i*8 +: 8];
		end
		
	endgenerate



endmodule 