module test_mem(input clk);


memory_mod(0,1,1,1,clk);




endmodule