module test_top(
	input clk,
	input sw1,
	input sw2,
	input sw3,
	output [7:0]leds
);
	//INSERE MATRIZ A 
	top(22'b10_11111111_00_000_000_0010, sw1, clk, leds);
	top(22'b10_11111111_00_000_010_0010, sw1, clk,  );
	top(22'b10_11111111_00_000_100_0010, sw1, clk,  );
	
	top(22'b10_11111111_00_001_001_0010, sw1, clk,  );
	top(22'b10_11111111_00_001_011_0010, sw1, clk,  );
	
	top(22'b10_11111111_00_010_000_0010, sw1, clk,  );
	top(22'b10_11111111_00_010_010_0010, sw1, clk,  );
	top(22'b10_11111111_00_010_100_0010, sw1, clk,  );

	top(22'b10_11111111_00_011_001_0010, sw1, clk,  );
	top(22'b10_11111111_00_011_011_0010, sw1, clk,  );
	
	top(22'b10_11111111_00_100_000_0010, sw1, clk,  );
	top(22'b10_11111111_00_100_010_0010, sw1, clk,  );
	top(22'b10_11111111_00_100_100_0010, sw1, clk,  );

	
	
	//INSERE MATRIZ B
	top(22'b10_11111111_01_000_000_0010, sw1, clk,  );
	top(22'b10_11111111_01_000_010_0010, sw1, clk,  );
	top(22'b10_11111111_01_000_100_0010, sw1, clk,  );
	
	top(22'b10_11111111_01_001_001_0010, sw1, clk,  );
	top(22'b10_11111111_01_001_011_0010, sw1, clk,  );
	
	top(22'b10_11111111_01_010_000_0010, sw1, clk,  );
	top(22'b10_11111111_01_010_010_0010, sw1, clk,  );
	top(22'b10_11111111_01_010_100_0010, sw1, clk,  );

	top(22'b10_11111111_01_011_001_0010, sw1, clk,  );
	top(22'b10_11111111_01_011_011_0010, sw1, clk,  );
	
	top(22'b10_11111111_01_100_000_0010, sw1, clk,  );
	top(22'b10_11111111_01_100_010_0010, sw1, clk,  );
	top(22'b10_11111111_01_100_100_0010, sw1, clk,  );
	
	
	//top(22'b00_00000000_00_000_000_0010, sw1, clk,  );
	
	
	
	
	
	
	
	
	
	
endmodule